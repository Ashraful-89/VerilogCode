module oRGate (a,b,sum);
input a ,b;
output sum;
or(sum,a,b);
endmodule
