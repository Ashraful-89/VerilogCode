module or_gate(a,b,sum);
	input a, b;
	output sum;
	or o1(sum, a, b);
endmodule
